`timescale 1ns / 1ps
module ext5(
    input [4:0]data_in,
    output [31:0]data_out
);
    assign data_out = {27'b0,data_in};

endmodule
